module segment(input [3:0] i, output reg [7:0] a, output reg [6:0] z);
always @(*)
case (i)
4'b0000 :  begin a=8'b11111110; z = 7'b1000000; end
4'b0001 :   begin a=8'b11111110; z = 7'b1111001; end
4'b0010 :   begin a=8'b11111110; z = 7'b0100100; end
4'b0011 :   begin a=8'b11111110; z = 7'b0110000; end
4'b0100 :  begin a=8'b11111110; z = 7'b0011001; end
4'b0101 :  begin a=8'b11111110; z = 7'b0010010; end
4'b0110 :  begin a=8'b11111110; z = 7'b0000010; end
4'b0111 :  begin a=8'b11111110; z = 7'b1111000; end
4'b1000 :   begin a=8'b11111110; z = 7'b0000000; end
4'b1001 :   begin a=8'b11111110; z = 7'b0010000; end
4'b1010 :   begin a=8'b11111110; z = 7'b0001000; end
4'b1011 :   begin a=8'b11111110; z = 7'b0000011; end
4'b1100 :  begin a=8'b11111110; z = 7'b1000110; end
4'b1101 :  begin a=8'b11111110; z = 7'b0100001; end
4'b1110 :  begin a=8'b11111110; z = 7'b0000110; end
4'b1111 :  begin a=8'b11111110; z = 7'b0001110; end
endcase    
endmodule
